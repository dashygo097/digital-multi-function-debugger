module sin_rom_a8d8(
	addr,
	clk, 
	q
);	

	parameter DATA_WIDTH=8;
	parameter ADDR_WIDTH=8;

	input clk;
	input [(ADDR_WIDTH-1):0] addr;
	output reg [(DATA_WIDTH-1):0] q;
	


	// Declare the ROM variable
	reg [DATA_WIDTH-1:0] rom[2**ADDR_WIDTH-1:0];

	initial begin
		rom[000] = 8'h7f; 
		rom[001] = 8'h82; 
		rom[002] = 8'h85; 
		rom[003] = 8'h88; 
		rom[004] = 8'h8b; 
		rom[005] = 8'h8f; 
		rom[006] = 8'h92; 
		rom[007] = 8'h95; 
		rom[008] = 8'h98; 
		rom[009] = 8'h9b; 
		rom[010] = 8'h9e; 
		rom[011] = 8'ha1; 
		rom[012] = 8'ha4; 
		rom[013] = 8'ha7; 
		rom[014] = 8'haa; 
		rom[015] = 8'had; 
		rom[016] = 8'hb0; 
		rom[017] = 8'hb2; 
		rom[018] = 8'hb5; 
		rom[019] = 8'hb8; 
		rom[020] = 8'hbb; 
		rom[021] = 8'hbe; 
		rom[022] = 8'hc0; 
		rom[023] = 8'hc3; 
		rom[024] = 8'hc6; 
		rom[025] = 8'hc8; 
		rom[026] = 8'hcb; 
		rom[027] = 8'hcd; 
		rom[028] = 8'hd0; 
		rom[029] = 8'hd2; 
		rom[030] = 8'hd4; 
		rom[031] = 8'hd7; 
		rom[032] = 8'hd9; 
		rom[033] = 8'hdb; 
		rom[034] = 8'hdd; 
		rom[035] = 8'hdf; 
		rom[036] = 8'he1; 
		rom[037] = 8'he3; 
		rom[038] = 8'he5; 
		rom[039] = 8'he7; 
		rom[040] = 8'he9; 
		rom[041] = 8'hea; 
		rom[042] = 8'hec; 
		rom[043] = 8'hee; 
		rom[044] = 8'hef; 
		rom[045] = 8'hf0; 
		rom[046] = 8'hf2; 
		rom[047] = 8'hf3; 
		rom[048] = 8'hf4; 
		rom[049] = 8'hf5; 
		rom[050] = 8'hf7; 
		rom[051] = 8'hf8; 
		rom[052] = 8'hf9; 
		rom[053] = 8'hf9; 
		rom[054] = 8'hfa; 
		rom[055] = 8'hfb; 
		rom[056] = 8'hfc; 
		rom[057] = 8'hfc; 
		rom[058] = 8'hfd; 
		rom[059] = 8'hfd; 
		rom[060] = 8'hfd; 
		rom[061] = 8'hfe; 
		rom[062] = 8'hfe; 
		rom[063] = 8'hfe; 
		rom[064] = 8'hfe; 
		rom[065] = 8'hfe; 
		rom[066] = 8'hfe; 
		rom[067] = 8'hfe; 
		rom[068] = 8'hfd; 
		rom[069] = 8'hfd; 
		rom[070] = 8'hfd; 
		rom[071] = 8'hfc; 
		rom[072] = 8'hfc; 
		rom[073] = 8'hfb; 
		rom[074] = 8'hfa; 
		rom[075] = 8'hf9; 
		rom[076] = 8'hf9; 
		rom[077] = 8'hf8; 
		rom[078] = 8'hf7; 
		rom[079] = 8'hf5; 
		rom[080] = 8'hf4; 
		rom[081] = 8'hf3; 
		rom[082] = 8'hf2; 
		rom[083] = 8'hf0; 
		rom[084] = 8'hef; 
		rom[085] = 8'hee; 
		rom[086] = 8'hec; 
		rom[087] = 8'hea; 
		rom[088] = 8'he9; 
		rom[089] = 8'he7; 
		rom[090] = 8'he5; 
		rom[091] = 8'he3; 
		rom[092] = 8'he1; 
		rom[093] = 8'hdf; 
		rom[094] = 8'hdd; 
		rom[095] = 8'hdb; 
		rom[096] = 8'hd9; 
		rom[097] = 8'hd7; 
		rom[098] = 8'hd4; 
		rom[099] = 8'hd2; 
		rom[100] = 8'hd0; 
		rom[101] = 8'hcd; 
		rom[102] = 8'hcb; 
		rom[103] = 8'hc8; 
		rom[104] = 8'hc6; 
		rom[105] = 8'hc3; 
		rom[106] = 8'hc0; 
		rom[107] = 8'hbe; 
		rom[108] = 8'hbb; 
		rom[109] = 8'hb8; 
		rom[110] = 8'hb5; 
		rom[111] = 8'hb2; 
		rom[112] = 8'hb0; 
		rom[113] = 8'had; 
		rom[114] = 8'haa; 
		rom[115] = 8'ha7; 
		rom[116] = 8'ha4; 
		rom[117] = 8'ha1; 
		rom[118] = 8'h9e; 
		rom[119] = 8'h9b; 
		rom[120] = 8'h98; 
		rom[121] = 8'h95; 
		rom[122] = 8'h92; 
		rom[123] = 8'h8f; 
		rom[124] = 8'h8b; 
		rom[125] = 8'h88; 
		rom[126] = 8'h85; 
		rom[127] = 8'h82; 
		rom[128] = 8'h7f; 
		rom[129] = 8'h7c; 
		rom[130] = 8'h79; 
		rom[131] = 8'h76; 
		rom[132] = 8'h73; 
		rom[133] = 8'h6f; 
		rom[134] = 8'h6c; 
		rom[135] = 8'h69; 
		rom[136] = 8'h66; 
		rom[137] = 8'h63; 
		rom[138] = 8'h60; 
		rom[139] = 8'h5d; 
		rom[140] = 8'h5a; 
		rom[141] = 8'h57; 
		rom[142] = 8'h54; 
		rom[143] = 8'h51; 
		rom[144] = 8'h4e; 
		rom[145] = 8'h4c; 
		rom[146] = 8'h49; 
		rom[147] = 8'h46; 
		rom[148] = 8'h43; 
		rom[149] = 8'h40; 
		rom[150] = 8'h3e; 
		rom[151] = 8'h3b; 
		rom[152] = 8'h38; 
		rom[153] = 8'h36; 
		rom[154] = 8'h33; 
		rom[155] = 8'h31; 
		rom[156] = 8'h2e; 
		rom[157] = 8'h2c; 
		rom[158] = 8'h2a; 
		rom[159] = 8'h27; 
		rom[160] = 8'h25; 
		rom[161] = 8'h23; 
		rom[162] = 8'h21; 
		rom[163] = 8'h1f; 
		rom[164] = 8'h1d; 
		rom[165] = 8'h1b; 
		rom[166] = 8'h19; 
		rom[167] = 8'h17; 
		rom[168] = 8'h15; 
		rom[169] = 8'h14; 
		rom[170] = 8'h12; 
		rom[171] = 8'h10; 
		rom[172] = 8'hf; 
		rom[173] = 8'he; 
		rom[174] = 8'hc; 
		rom[175] = 8'hb; 
		rom[176] = 8'ha; 
		rom[177] = 8'h9; 
		rom[178] = 8'h7; 
		rom[179] = 8'h6; 
		rom[180] = 8'h5; 
		rom[181] = 8'h5; 
		rom[182] = 8'h4; 
		rom[183] = 8'h3; 
		rom[184] = 8'h2; 
		rom[185] = 8'h2; 
		rom[186] = 8'h1; 
		rom[187] = 8'h1; 
		rom[188] = 8'h1; 
		rom[189] = 8'h0; 
		rom[190] = 8'h0; 
		rom[191] = 8'h0; 
		rom[192] = 8'h0; 
		rom[193] = 8'h0; 
		rom[194] = 8'h0; 
		rom[195] = 8'h0; 
		rom[196] = 8'h1; 
		rom[197] = 8'h1; 
		rom[198] = 8'h1; 
		rom[199] = 8'h2; 
		rom[200] = 8'h2; 
		rom[201] = 8'h3; 
		rom[202] = 8'h4; 
		rom[203] = 8'h5; 
		rom[204] = 8'h5; 
		rom[205] = 8'h6; 
		rom[206] = 8'h7; 
		rom[207] = 8'h9; 
		rom[208] = 8'ha; 
		rom[209] = 8'hb; 
		rom[210] = 8'hc; 
		rom[211] = 8'he; 
		rom[212] = 8'hf; 
		rom[213] = 8'h10; 
		rom[214] = 8'h12; 
		rom[215] = 8'h14; 
		rom[216] = 8'h15; 
		rom[217] = 8'h17; 
		rom[218] = 8'h19; 
		rom[219] = 8'h1b; 
		rom[220] = 8'h1d; 
		rom[221] = 8'h1f; 
		rom[222] = 8'h21; 
		rom[223] = 8'h23; 
		rom[224] = 8'h25; 
		rom[225] = 8'h27; 
		rom[226] = 8'h2a; 
		rom[227] = 8'h2c; 
		rom[228] = 8'h2e; 
		rom[229] = 8'h31; 
		rom[230] = 8'h33; 
		rom[231] = 8'h36; 
		rom[232] = 8'h38; 
		rom[233] = 8'h3b; 
		rom[234] = 8'h3e; 
		rom[235] = 8'h40; 
		rom[236] = 8'h43; 
		rom[237] = 8'h46; 
		rom[238] = 8'h49; 
		rom[239] = 8'h4c; 
		rom[240] = 8'h4e; 
		rom[241] = 8'h51; 
		rom[242] = 8'h54; 
		rom[243] = 8'h57; 
		rom[244] = 8'h5a; 
		rom[245] = 8'h5d; 
		rom[246] = 8'h60; 
		rom[247] = 8'h63; 
		rom[248] = 8'h66; 
		rom[249] = 8'h69; 
		rom[250] = 8'h6c; 
		rom[251] = 8'h6f; 
		rom[252] = 8'h73; 
		rom[253] = 8'h76; 
		rom[254] = 8'h79; 
		rom[255] = 8'h7c;
	end

	always @ (posedge clk)
	begin
		q <= rom[addr];
	end

endmodule
