//Copyright (C)2014-2023 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.9 Beta-3
//Part Number: GW5A-LV25UG324ES
//Device: GW5A-25
//Device Version: A
//Created Time: Wed Sep 13 11:40:51 2023

module rom_triangular (dout, clk, oce, ce, reset, ad);

output [13:0] dout;
input clk;
input oce;
input ce;
input reset;
input [11:0] ad;

wire [27:0] prom_inst_0_dout_w;
wire [27:0] prom_inst_1_dout_w;
wire [27:0] prom_inst_2_dout_w;
wire [29:0] prom_inst_3_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[27:0],dout[3:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 4;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h8080808080808080808080808080808080808080808080808080808080808080;
defparam prom_inst_0.INIT_RAM_01 = 256'h8080808080808080808080808080808080808080808080808080808080808080;
defparam prom_inst_0.INIT_RAM_02 = 256'h8080808080808080808080808080808080808080808080808080808080808080;
defparam prom_inst_0.INIT_RAM_03 = 256'h8080808080808080808080808080808080808080808080808080808080808080;
defparam prom_inst_0.INIT_RAM_04 = 256'h8080808080808080808080808080808080808080808080808080808080808080;
defparam prom_inst_0.INIT_RAM_05 = 256'h8080808080808080808080808080808080808080808080808080808080808080;
defparam prom_inst_0.INIT_RAM_06 = 256'h8080808080808080808080808080808080808080808080808080808080808080;
defparam prom_inst_0.INIT_RAM_07 = 256'h8080808080808080808080808080808080808080808080808080808080808080;
defparam prom_inst_0.INIT_RAM_08 = 256'h8080808080808080808080808080808080808080808080808080808080808080;
defparam prom_inst_0.INIT_RAM_09 = 256'h8080808080808080808080808080808080808080808080808080808080808080;
defparam prom_inst_0.INIT_RAM_0A = 256'h8080808080808080808080808080808080808080808080808080808080808080;
defparam prom_inst_0.INIT_RAM_0B = 256'h8080808080808080808080808080808080808080808080808080808080808080;
defparam prom_inst_0.INIT_RAM_0C = 256'h8080808080808080808080808080808080808080808080808080808080808080;
defparam prom_inst_0.INIT_RAM_0D = 256'h8080808080808080808080808080808080808080808080808080808080808080;
defparam prom_inst_0.INIT_RAM_0E = 256'h8080808080808080808080808080808080808080808080808080808080808080;
defparam prom_inst_0.INIT_RAM_0F = 256'h8080808080808080808080808080808080808080808080808080808080808080;
defparam prom_inst_0.INIT_RAM_10 = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F70;
defparam prom_inst_0.INIT_RAM_11 = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_0.INIT_RAM_12 = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_0.INIT_RAM_13 = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_0.INIT_RAM_14 = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_0.INIT_RAM_15 = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_0.INIT_RAM_16 = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_0.INIT_RAM_17 = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_0.INIT_RAM_18 = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_0.INIT_RAM_19 = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_0.INIT_RAM_1A = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_0.INIT_RAM_1B = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_0.INIT_RAM_1C = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_0.INIT_RAM_1D = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_0.INIT_RAM_1E = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_0.INIT_RAM_1F = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_0.INIT_RAM_20 = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_0.INIT_RAM_21 = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_0.INIT_RAM_22 = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_0.INIT_RAM_23 = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_0.INIT_RAM_24 = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_0.INIT_RAM_25 = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_0.INIT_RAM_26 = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_0.INIT_RAM_27 = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_0.INIT_RAM_28 = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_0.INIT_RAM_29 = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_0.INIT_RAM_2A = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_0.INIT_RAM_2B = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_0.INIT_RAM_2C = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_0.INIT_RAM_2D = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_0.INIT_RAM_2E = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_0.INIT_RAM_2F = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_0.INIT_RAM_30 = 256'h8080808080808080808080808080808080808080808080808080808080808080;
defparam prom_inst_0.INIT_RAM_31 = 256'h8080808080808080808080808080808080808080808080808080808080808080;
defparam prom_inst_0.INIT_RAM_32 = 256'h8080808080808080808080808080808080808080808080808080808080808080;
defparam prom_inst_0.INIT_RAM_33 = 256'h8080808080808080808080808080808080808080808080808080808080808080;
defparam prom_inst_0.INIT_RAM_34 = 256'h8080808080808080808080808080808080808080808080808080808080808080;
defparam prom_inst_0.INIT_RAM_35 = 256'h8080808080808080808080808080808080808080808080808080808080808080;
defparam prom_inst_0.INIT_RAM_36 = 256'h8080808080808080808080808080808080808080808080808080808080808080;
defparam prom_inst_0.INIT_RAM_37 = 256'h8080808080808080808080808080808080808080808080808080808080808080;
defparam prom_inst_0.INIT_RAM_38 = 256'h8080808080808080808080808080808080808080808080808080808080808080;
defparam prom_inst_0.INIT_RAM_39 = 256'h8080808080808080808080808080808080808080808080808080808080808080;
defparam prom_inst_0.INIT_RAM_3A = 256'h8080808080808080808080808080808080808080808080808080808080808080;
defparam prom_inst_0.INIT_RAM_3B = 256'h8080808080808080808080808080808080808080808080808080808080808080;
defparam prom_inst_0.INIT_RAM_3C = 256'h8080808080808080808080808080808080808080808080808080808080808080;
defparam prom_inst_0.INIT_RAM_3D = 256'h8080808080808080808080808080808080808080808080808080808080808080;
defparam prom_inst_0.INIT_RAM_3E = 256'h8080808080808080808080808080808080808080808080808080808080808080;
defparam prom_inst_0.INIT_RAM_3F = 256'h8080808080808080808080808080808080808080808080808080808080808080;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[27:0],dout[7:4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 4;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'hFFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100;
defparam prom_inst_1.INIT_RAM_01 = 256'hFFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100;
defparam prom_inst_1.INIT_RAM_02 = 256'hFFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100;
defparam prom_inst_1.INIT_RAM_03 = 256'hFFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100;
defparam prom_inst_1.INIT_RAM_04 = 256'hFFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100;
defparam prom_inst_1.INIT_RAM_05 = 256'hFFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100;
defparam prom_inst_1.INIT_RAM_06 = 256'hFFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100;
defparam prom_inst_1.INIT_RAM_07 = 256'hFFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100;
defparam prom_inst_1.INIT_RAM_08 = 256'hFFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100;
defparam prom_inst_1.INIT_RAM_09 = 256'hFFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100;
defparam prom_inst_1.INIT_RAM_0A = 256'hFFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100;
defparam prom_inst_1.INIT_RAM_0B = 256'hFFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100;
defparam prom_inst_1.INIT_RAM_0C = 256'hFFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100;
defparam prom_inst_1.INIT_RAM_0D = 256'hFFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100;
defparam prom_inst_1.INIT_RAM_0E = 256'hFFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100;
defparam prom_inst_1.INIT_RAM_0F = 256'hFFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100;
defparam prom_inst_1.INIT_RAM_10 = 256'hFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA998877665544332211000;
defparam prom_inst_1.INIT_RAM_11 = 256'hFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100F;
defparam prom_inst_1.INIT_RAM_12 = 256'hFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100F;
defparam prom_inst_1.INIT_RAM_13 = 256'hFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100F;
defparam prom_inst_1.INIT_RAM_14 = 256'hFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100F;
defparam prom_inst_1.INIT_RAM_15 = 256'hFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100F;
defparam prom_inst_1.INIT_RAM_16 = 256'hFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100F;
defparam prom_inst_1.INIT_RAM_17 = 256'hFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100F;
defparam prom_inst_1.INIT_RAM_18 = 256'hFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100F;
defparam prom_inst_1.INIT_RAM_19 = 256'hFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100F;
defparam prom_inst_1.INIT_RAM_1A = 256'hFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100F;
defparam prom_inst_1.INIT_RAM_1B = 256'hFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100F;
defparam prom_inst_1.INIT_RAM_1C = 256'hFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100F;
defparam prom_inst_1.INIT_RAM_1D = 256'hFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100F;
defparam prom_inst_1.INIT_RAM_1E = 256'hFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100F;
defparam prom_inst_1.INIT_RAM_1F = 256'hFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100F;
defparam prom_inst_1.INIT_RAM_20 = 256'h00112233445566778899AABBCCDDEEFF00112233445566778899AABBCCDDEEFF;
defparam prom_inst_1.INIT_RAM_21 = 256'h00112233445566778899AABBCCDDEEFF00112233445566778899AABBCCDDEEFF;
defparam prom_inst_1.INIT_RAM_22 = 256'h00112233445566778899AABBCCDDEEFF00112233445566778899AABBCCDDEEFF;
defparam prom_inst_1.INIT_RAM_23 = 256'h00112233445566778899AABBCCDDEEFF00112233445566778899AABBCCDDEEFF;
defparam prom_inst_1.INIT_RAM_24 = 256'h00112233445566778899AABBCCDDEEFF00112233445566778899AABBCCDDEEFF;
defparam prom_inst_1.INIT_RAM_25 = 256'h00112233445566778899AABBCCDDEEFF00112233445566778899AABBCCDDEEFF;
defparam prom_inst_1.INIT_RAM_26 = 256'h00112233445566778899AABBCCDDEEFF00112233445566778899AABBCCDDEEFF;
defparam prom_inst_1.INIT_RAM_27 = 256'h00112233445566778899AABBCCDDEEFF00112233445566778899AABBCCDDEEFF;
defparam prom_inst_1.INIT_RAM_28 = 256'h00112233445566778899AABBCCDDEEFF00112233445566778899AABBCCDDEEFF;
defparam prom_inst_1.INIT_RAM_29 = 256'h00112233445566778899AABBCCDDEEFF00112233445566778899AABBCCDDEEFF;
defparam prom_inst_1.INIT_RAM_2A = 256'h00112233445566778899AABBCCDDEEFF00112233445566778899AABBCCDDEEFF;
defparam prom_inst_1.INIT_RAM_2B = 256'h00112233445566778899AABBCCDDEEFF00112233445566778899AABBCCDDEEFF;
defparam prom_inst_1.INIT_RAM_2C = 256'h00112233445566778899AABBCCDDEEFF00112233445566778899AABBCCDDEEFF;
defparam prom_inst_1.INIT_RAM_2D = 256'h00112233445566778899AABBCCDDEEFF00112233445566778899AABBCCDDEEFF;
defparam prom_inst_1.INIT_RAM_2E = 256'h00112233445566778899AABBCCDDEEFF00112233445566778899AABBCCDDEEFF;
defparam prom_inst_1.INIT_RAM_2F = 256'h00112233445566778899AABBCCDDEEFF00112233445566778899AABBCCDDEEFF;
defparam prom_inst_1.INIT_RAM_30 = 256'h0112233445566778899AABBCCDDEEFF00112233445566778899AABBCCDDEEFF0;
defparam prom_inst_1.INIT_RAM_31 = 256'h0112233445566778899AABBCCDDEEFF00112233445566778899AABBCCDDEEFF0;
defparam prom_inst_1.INIT_RAM_32 = 256'h0112233445566778899AABBCCDDEEFF00112233445566778899AABBCCDDEEFF0;
defparam prom_inst_1.INIT_RAM_33 = 256'h0112233445566778899AABBCCDDEEFF00112233445566778899AABBCCDDEEFF0;
defparam prom_inst_1.INIT_RAM_34 = 256'h0112233445566778899AABBCCDDEEFF00112233445566778899AABBCCDDEEFF0;
defparam prom_inst_1.INIT_RAM_35 = 256'h0112233445566778899AABBCCDDEEFF00112233445566778899AABBCCDDEEFF0;
defparam prom_inst_1.INIT_RAM_36 = 256'h0112233445566778899AABBCCDDEEFF00112233445566778899AABBCCDDEEFF0;
defparam prom_inst_1.INIT_RAM_37 = 256'h0112233445566778899AABBCCDDEEFF00112233445566778899AABBCCDDEEFF0;
defparam prom_inst_1.INIT_RAM_38 = 256'h0112233445566778899AABBCCDDEEFF00112233445566778899AABBCCDDEEFF0;
defparam prom_inst_1.INIT_RAM_39 = 256'h0112233445566778899AABBCCDDEEFF00112233445566778899AABBCCDDEEFF0;
defparam prom_inst_1.INIT_RAM_3A = 256'h0112233445566778899AABBCCDDEEFF00112233445566778899AABBCCDDEEFF0;
defparam prom_inst_1.INIT_RAM_3B = 256'h0112233445566778899AABBCCDDEEFF00112233445566778899AABBCCDDEEFF0;
defparam prom_inst_1.INIT_RAM_3C = 256'h0112233445566778899AABBCCDDEEFF00112233445566778899AABBCCDDEEFF0;
defparam prom_inst_1.INIT_RAM_3D = 256'h0112233445566778899AABBCCDDEEFF00112233445566778899AABBCCDDEEFF0;
defparam prom_inst_1.INIT_RAM_3E = 256'h0112233445566778899AABBCCDDEEFF00112233445566778899AABBCCDDEEFF0;
defparam prom_inst_1.INIT_RAM_3F = 256'h0112233445566778899AABBCCDDEEFF00112233445566778899AABBCCDDEEFF0;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[27:0],dout[11:8]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 4;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'h1111111111111111111111111111111100000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_01 = 256'h3333333333333333333333333333333322222222222222222222222222222222;
defparam prom_inst_2.INIT_RAM_02 = 256'h5555555555555555555555555555555544444444444444444444444444444444;
defparam prom_inst_2.INIT_RAM_03 = 256'h7777777777777777777777777777777766666666666666666666666666666666;
defparam prom_inst_2.INIT_RAM_04 = 256'h9999999999999999999999999999999988888888888888888888888888888888;
defparam prom_inst_2.INIT_RAM_05 = 256'hBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_2.INIT_RAM_06 = 256'hDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCC;
defparam prom_inst_2.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam prom_inst_2.INIT_RAM_08 = 256'h1111111111111111111111111111111100000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_09 = 256'h3333333333333333333333333333333322222222222222222222222222222222;
defparam prom_inst_2.INIT_RAM_0A = 256'h5555555555555555555555555555555544444444444444444444444444444444;
defparam prom_inst_2.INIT_RAM_0B = 256'h7777777777777777777777777777777766666666666666666666666666666666;
defparam prom_inst_2.INIT_RAM_0C = 256'h9999999999999999999999999999999988888888888888888888888888888888;
defparam prom_inst_2.INIT_RAM_0D = 256'hBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_2.INIT_RAM_0E = 256'hDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCC;
defparam prom_inst_2.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam prom_inst_2.INIT_RAM_10 = 256'h1111111111111111111111111111111000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_11 = 256'h3333333333333333333333333333333222222222222222222222222222222221;
defparam prom_inst_2.INIT_RAM_12 = 256'h5555555555555555555555555555555444444444444444444444444444444443;
defparam prom_inst_2.INIT_RAM_13 = 256'h7777777777777777777777777777777666666666666666666666666666666665;
defparam prom_inst_2.INIT_RAM_14 = 256'h9999999999999999999999999999999888888888888888888888888888888887;
defparam prom_inst_2.INIT_RAM_15 = 256'hBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9;
defparam prom_inst_2.INIT_RAM_16 = 256'hDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCB;
defparam prom_inst_2.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEED;
defparam prom_inst_2.INIT_RAM_18 = 256'h111111111111111111111111111111100000000000000000000000000000000F;
defparam prom_inst_2.INIT_RAM_19 = 256'h3333333333333333333333333333333222222222222222222222222222222221;
defparam prom_inst_2.INIT_RAM_1A = 256'h5555555555555555555555555555555444444444444444444444444444444443;
defparam prom_inst_2.INIT_RAM_1B = 256'h7777777777777777777777777777777666666666666666666666666666666665;
defparam prom_inst_2.INIT_RAM_1C = 256'h9999999999999999999999999999999888888888888888888888888888888887;
defparam prom_inst_2.INIT_RAM_1D = 256'hBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9;
defparam prom_inst_2.INIT_RAM_1E = 256'hDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCB;
defparam prom_inst_2.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEED;
defparam prom_inst_2.INIT_RAM_20 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_21 = 256'hCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD;
defparam prom_inst_2.INIT_RAM_22 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB;
defparam prom_inst_2.INIT_RAM_23 = 256'h8888888888888888888888888888888899999999999999999999999999999999;
defparam prom_inst_2.INIT_RAM_24 = 256'h6666666666666666666666666666666677777777777777777777777777777777;
defparam prom_inst_2.INIT_RAM_25 = 256'h4444444444444444444444444444444455555555555555555555555555555555;
defparam prom_inst_2.INIT_RAM_26 = 256'h2222222222222222222222222222222233333333333333333333333333333333;
defparam prom_inst_2.INIT_RAM_27 = 256'h0000000000000000000000000000000011111111111111111111111111111111;
defparam prom_inst_2.INIT_RAM_28 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_29 = 256'hCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD;
defparam prom_inst_2.INIT_RAM_2A = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB;
defparam prom_inst_2.INIT_RAM_2B = 256'h8888888888888888888888888888888899999999999999999999999999999999;
defparam prom_inst_2.INIT_RAM_2C = 256'h6666666666666666666666666666666677777777777777777777777777777777;
defparam prom_inst_2.INIT_RAM_2D = 256'h4444444444444444444444444444444455555555555555555555555555555555;
defparam prom_inst_2.INIT_RAM_2E = 256'h2222222222222222222222222222222233333333333333333333333333333333;
defparam prom_inst_2.INIT_RAM_2F = 256'h0000000000000000000000000000000011111111111111111111111111111111;
defparam prom_inst_2.INIT_RAM_30 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0;
defparam prom_inst_2.INIT_RAM_31 = 256'hCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDE;
defparam prom_inst_2.INIT_RAM_32 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBC;
defparam prom_inst_2.INIT_RAM_33 = 256'h888888888888888888888888888888899999999999999999999999999999999A;
defparam prom_inst_2.INIT_RAM_34 = 256'h6666666666666666666666666666666777777777777777777777777777777778;
defparam prom_inst_2.INIT_RAM_35 = 256'h4444444444444444444444444444444555555555555555555555555555555556;
defparam prom_inst_2.INIT_RAM_36 = 256'h2222222222222222222222222222222333333333333333333333333333333334;
defparam prom_inst_2.INIT_RAM_37 = 256'h0000000000000000000000000000000111111111111111111111111111111112;
defparam prom_inst_2.INIT_RAM_38 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0;
defparam prom_inst_2.INIT_RAM_39 = 256'hCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDE;
defparam prom_inst_2.INIT_RAM_3A = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBC;
defparam prom_inst_2.INIT_RAM_3B = 256'h888888888888888888888888888888899999999999999999999999999999999A;
defparam prom_inst_2.INIT_RAM_3C = 256'h6666666666666666666666666666666777777777777777777777777777777778;
defparam prom_inst_2.INIT_RAM_3D = 256'h4444444444444444444444444444444555555555555555555555555555555556;
defparam prom_inst_2.INIT_RAM_3E = 256'h2222222222222222222222222222222333333333333333333333333333333334;
defparam prom_inst_2.INIT_RAM_3F = 256'h0000000000000000000000000000000111111111111111111111111111111112;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[29:0],dout[13:12]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({gw_gnd,ad[11:0],gw_gnd})
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 2;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_04 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
defparam prom_inst_3.INIT_RAM_05 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
defparam prom_inst_3.INIT_RAM_06 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
defparam prom_inst_3.INIT_RAM_07 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
defparam prom_inst_3.INIT_RAM_08 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_3.INIT_RAM_09 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_3.INIT_RAM_0A = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_3.INIT_RAM_0B = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_3.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE;
defparam prom_inst_3.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_14 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_3.INIT_RAM_15 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_3.INIT_RAM_16 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_3.INIT_RAM_17 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_3.INIT_RAM_18 = 256'h5555555555555555555555555555555555555555555555555555555555555556;
defparam prom_inst_3.INIT_RAM_19 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
defparam prom_inst_3.INIT_RAM_1A = 256'h5555555555555555555555555555555555555555555555555555555555555555;
defparam prom_inst_3.INIT_RAM_1B = 256'h5555555555555555555555555555555555555555555555555555555555555555;
defparam prom_inst_3.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_3.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule //rom_triangular
