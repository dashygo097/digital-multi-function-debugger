//Copyright (C)2014-2023 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.9 Beta-3
//Part Number: GW5A-LV25UG324ES
//Device: GW5A-25
//Device Version: A
//Created Time: Fri Sep 08 14:47:18 2023

module rom_sine (dout, clk, oce, ce, reset, ad);

output [13:0] dout;
input clk;
input oce;
input ce;
input reset;
input [11:0] ad;

wire [27:0] prom_inst_0_dout_w;
wire [27:0] prom_inst_1_dout_w;
wire [27:0] prom_inst_2_dout_w;
wire [29:0] prom_inst_3_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[27:0],dout[3:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 4;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h59C037AE158CF36AD147BE259C037AD148BF269C037AE158BF269D047AE158CF;
defparam prom_inst_0.INIT_RAM_01 = 256'h148CF37AE259C047BF269D148BF36AD148CF36AD148CF36AD148BF269D047BE2;
defparam prom_inst_0.INIT_RAM_02 = 256'hD159D048C048C048CF37BF37AE26AE159D148C047BF36AE259D148CF37BE269D;
defparam prom_inst_0.INIT_RAM_03 = 256'h26BF38C059D26AF37B048C159D26AE26BF37BF38C048C048C059D159D159D159;
defparam prom_inst_0.INIT_RAM_04 = 256'h9E38D26B05AF38D27B05AE38C16AF48D26B049D27B049D26BF48D16AF38C059E;
defparam prom_inst_0.INIT_RAM_05 = 256'hB16C17C27D28D28D38D38D38D28D28D27C27C16B16B05AF49E39E38D27C05AF4;
defparam prom_inst_0.INIT_RAM_06 = 256'h28E4B17D3A06C28E4B17D39F5B17D38E4A06C27D39F4A06B17D28E39F4AF5B06;
defparam prom_inst_0.INIT_RAM_07 = 256'h6D4B2907E5C3A18F6D4B18F6D3A18E5C2906D4A17E5B28F5C29F5C29F5C28F5B;
defparam prom_inst_0.INIT_RAM_08 = 256'h3B3B3B3A2A2A2A19191808F7F7E6D5D4C3B2A1908F6E5D4B3A1907E6D4B2A18F;
defparam prom_inst_0.INIT_RAM_09 = 256'h3C5E6F81A3C5D6F8192B3C5D6F7081A2B3C4C5D6E6F7F80819192A2A2A2A3B3B;
defparam prom_inst_0.INIT_RAM_0A = 256'h1B5F93D71B5F82C6093D70A4D71A4E71A4D70A3C6F92B5E70A3C5F81A3C5E71A;
defparam prom_inst_0.INIT_RAM_0B = 256'hA50B61C73E94E94FA50B60B61B61C61C61B60B60B5FA4F93E82D71B60A4E93D7;
defparam prom_inst_0.INIT_RAM_0C = 256'hA62FB730C840C851D951D950C840C83FB72EA51D840B72E950B72E940B62D83E;
defparam prom_inst_0.INIT_RAM_0D = 256'hEC9742FCA752FCA741FC9630DB852FC952FC9630C963FC952FB841DA63FC851D;
defparam prom_inst_0.INIT_RAM_0E = 256'h54310FDCB9865320FDCA875320EDB975320ECA86420ECA8531FDA8641FDA8531;
defparam prom_inst_0.INIT_RAM_0F = 256'hEEEEEEEDDDDDCCCCBBBAA99887766554432210FFEDCBAA9876543210FECBA987;
defparam prom_inst_0.INIT_RAM_10 = 256'h89ABCEF0123456789AABCDEFF01223445566778899AABBBCCCCDDDDDEEEEEEEE;
defparam prom_inst_0.INIT_RAM_11 = 256'h358ADF1468ADF1358ACE02468ACE023579BDE023578ACDF0235689BCDF013457;
defparam prom_inst_0.INIT_RAM_12 = 256'h158CF36AD148BF259CF369C0369CF259CF258BD0369CF147ACF257ACF2479CE1;
defparam prom_inst_0.INIT_RAM_13 = 256'h38D26B049E27B059E27B048D15AE27BF38C048C059D159D158C048C037BF26AD;
defparam prom_inst_0.INIT_RAM_14 = 256'hD39E4A06B17D28E39F4AF5B06B06B16C16C16B16B06B05AF49E49E37C16B05AE;
defparam prom_inst_0.INIT_RAM_15 = 256'h17E5C3A18F5C3A07E5B29F6C3A07D4A17E4A17D4A07D3906C28F5B17D39F5B17;
defparam prom_inst_0.INIT_RAM_16 = 256'h3B3A2A2A2A29191808F7F6E6D5C4C3B2A1807F6D5C3B2918F6D5C3A18F6E5C3A;
defparam prom_inst_0.INIT_RAM_17 = 256'h81A2B4D6E7091A3B4D5E6F8091A2B3C4D5D6E7F7F80819191A2A2A2A3B3B3B3B;
defparam prom_inst_0.INIT_RAM_18 = 256'h5F82C5F92C5F92C5F82B5E71A4D6092C5E81A3D6F81B4D6F81A3C5E7092B4D6F;
defparam prom_inst_0.INIT_RAM_19 = 256'h0B5FA4F93E82D71B60A4F93D72C60A4E83D71B5F93D71B4E82C60A3D71B4E82B;
defparam prom_inst_0.INIT_RAM_1A = 256'hFA50C72D83E93E94FA50B61B61C72C72D82D82D83D83D83D82D82D72C71C61B6;
defparam prom_inst_0.INIT_RAM_1B = 256'h950C83FA61D84FB62D940B72D940B62D84FA61C83EA50B72D83FA50B62D83E94;
defparam prom_inst_0.INIT_RAM_1C = 256'h51D951D951D950C840C840C83FB73FB62EA62D951C840B73FA62D950C83FB62E;
defparam prom_inst_0.INIT_RAM_1D = 256'h962EB73FC841D952EA63FB740C841D951EA62EA73FB73FC840C840C840D951D9;
defparam prom_inst_0.INIT_RAM_1E = 256'hEB740D962FB841DA63FC841DA63FC841DA63FB841D962FB740C952EA73FC841D;
defparam prom_inst_0.INIT_RAM_1F = 256'hC851EA740D962FB851EA730C962FB841DA730C952EB741DA63FC851EA730C952;
defparam prom_inst_0.INIT_RAM_20 = 256'h952EB740D962FB841DA730C952EB741DA63FC852EB740D963FC851EA740D962F;
defparam prom_inst_0.INIT_RAM_21 = 256'hDA62FB740C952EA73FC851DA63FB841DA62FB841DA62FB841DA63FC851EA730C;
defparam prom_inst_0.INIT_RAM_22 = 256'h1D951EA62EA62EA62FB73FB740C840D951DA62EA73FB840C951DA62FB730C851;
defparam prom_inst_0.INIT_RAM_23 = 256'hC83FB62E951C84FB73EA62D951C840C83FB73FB62EA62EA62E951D951D951D95;
defparam prom_inst_0.INIT_RAM_24 = 256'h50B61C83E94FB61C73E940B62D84FA61C83EA51C73EA51C83FA61D84FB62E950;
defparam prom_inst_0.INIT_RAM_25 = 256'h3D82D72C71C61C61B61B61B61C61C61C72C72D83D83E94FA50B50B61C72E94FA;
defparam prom_inst_0.INIT_RAM_26 = 256'hC60A3D71B4E82C60A3D71B5F93D71B60A4E82C71B5FA4E83D71C60B5FA4F93E8;
defparam prom_inst_0.INIT_RAM_27 = 256'h81A3C5E7092B4D6F81A3D6F81B4D6092C5E81A4D7093C6F92C5F92C5F92C6F93;
defparam prom_inst_0.INIT_RAM_28 = 256'hB3B3B3B4C4C4C4D5D5D6E6F7F708191A2B3C4D5E6F8091A3B4D5E7081A3C4D6F;
defparam prom_inst_0.INIT_RAM_29 = 256'hB2908F6D4B2918F6D5C3B2918F7E6D4C3B2A291808F7F6E6D5D5C4C4C4C4B3B3;
defparam prom_inst_0.INIT_RAM_2A = 256'hD39F5B17D39F6C28E5B17E4A17D4A07D4A17E4B28F5C3907E4B29F6D4B2907D4;
defparam prom_inst_0.INIT_RAM_2B = 256'h49E38D27B05A05AF49E38E38D38D28D28D38E38E39F4AF5B06C17D38E4A05B17;
defparam prom_inst_0.INIT_RAM_2C = 256'h48CF37BE26AE269D159D159E26AE26BF37C049D16AE37C059E37C05AE38C16B0;
defparam prom_inst_0.INIT_RAM_2D = 256'h0257ACF2479CF247ADF258BE1369CF259CF258BE258BF259CF36AD148BF269D1;
defparam prom_inst_0.INIT_RAM_2E = 256'h9ABDEF1235689BCEF124679BCE013579BCE02468ACE02469BDF1468ADF1469BD;
defparam prom_inst_0.INIT_RAM_2F = 256'h0000000111112222333445566778899AABCCDEFF01234456789ABCDEF0234567;
defparam prom_inst_0.INIT_RAM_30 = 256'h654320FEDCBA98765443210FFEDCCBAA99887766554433322221111100000000;
defparam prom_inst_0.INIT_RAM_31 = 256'hB9641FDA8641FDB96420ECA86420ECB975310ECB976421FECB9865321FEDBA97;
defparam prom_inst_0.INIT_RAM_32 = 256'hD962FB841DA63FC952FB852EB852FC952FC9631EB852FDA742FC9742FCA7520D;
defparam prom_inst_0.INIT_RAM_33 = 256'hB61C83EA50C73E950C73EA61D940C73FB62EA62E951D951D962EA62EB73FC841;
defparam prom_inst_0.INIT_RAM_34 = 256'h1B50A4E83D71C60B5FA4F93E83E83D82D82D83D83E83E94FA50A50B72D83E940;
defparam prom_inst_0.INIT_RAM_35 = 256'hD7092B4D6F92B4E7093C5F82B4E71A4D70A4D71A4E71B5E82C6F93D71B5F93D7;
defparam prom_inst_0.INIT_RAM_36 = 256'hB3B4C4C4C4C5D5D6E6F7F808192A2B3C4D6E7F8192B3C5D6F8192B4D6F8092B4;
defparam prom_inst_0.INIT_RAM_37 = 256'h6D4C3A1807E5D4B3A1908F6E5D4C3B2A191807F7F6E6D5D5D4C4C4C4B3B3B3B3;
defparam prom_inst_0.INIT_RAM_38 = 256'h9F6C29F5C29F5C29F6C3907D4A18E5C2906D4B18F6D3A18F6D4B2907E5C3A18F;
defparam prom_inst_0.INIT_RAM_39 = 256'hE39F4AF5B06C17D38E4AF5B17C28E4A06B17D39F5B17D3A06C28E4B17D3A06C3;
defparam prom_inst_0.INIT_RAM_3A = 256'hF49E27C16B05B05AF49E38D38D27C27C16C16C16B16B16B16C16C17C27D28D38;
defparam prom_inst_0.INIT_RAM_3B = 256'h59E26BF48D16AF38C15AE37C15AE38C16AF48D26B049E37C16BF49E38C16B05A;
defparam prom_inst_0.INIT_RAM_3C = 256'h9D159D159D159E26AE26AE26BF37BF38C048C159D26AE37BF48C159E26BF38C0;
defparam prom_inst_0.INIT_RAM_3D = 256'h58C037BF26AD159C048BF37AE26AD159D048C047BF37BF26AE26AE26AE159D15;
defparam prom_inst_0.INIT_RAM_3E = 256'h037AE158CF36AD148BF26AD148BF26AD148BF36AD158CF37AE259C047BF26AD1;
defparam prom_inst_0.INIT_RAM_3F = 256'h269D047AE158CF369D047BE258CF36AD147BE259C037AD148BF269D047BE259C;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[27:0],dout[7:4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 4;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'h10FFEDCBBA9877654432100FEDDCBA9987655432210FEEDCBAA987765433210F;
defparam prom_inst_1.INIT_RAM_01 = 256'h3210FFEDCCBA9987655432210FEEDCBBA9877654432100FEDDCBA99876654322;
defparam prom_inst_1.INIT_RAM_02 = 256'h332100FEDDCBAA9876654332100FEDDCBAA9877654332100FEDDCBA998766543;
defparam prom_inst_1.INIT_RAM_03 = 256'h32100FEEDCBBA98876654332100FEDDCBAA9877655432210FFEDCCBA99876654;
defparam prom_inst_1.INIT_RAM_04 = 256'h0FFEDDCBBA98876654432110FFEDCCBAA98876554332100FEDDCBBA988766543;
defparam prom_inst_1.INIT_RAM_05 = 256'hBBA998776554332110FFEDDCBBA998776554332110FFEDCCBAA9887665443211;
defparam prom_inst_1.INIT_RAM_06 = 256'h4322110FFEEDCCBAA9987765544322100FFEDDCBBA9988766544322100FEEDDC;
defparam prom_inst_1.INIT_RAM_07 = 256'h98877665443322100FFEEDCCBBAA98877665443321100FEEDDCBBAA988776554;
defparam prom_inst_1.INIT_RAM_08 = 256'hBAA9988776655443322110FFEEDDCCBBAA9988776554433221100FEEDDCCBBA9;
defparam prom_inst_1.INIT_RAM_09 = 256'h988776665544332221100FFEEDDDCCBBAA998877665544433221100FFEEDDCCB;
defparam prom_inst_1.INIT_RAM_0A = 256'h322111000FFEEEDDDCCBBBAA9998877766555443322211000FFEEDDDCCBBAAA9;
defparam prom_inst_1.INIT_RAM_0B = 256'h8887776665554443333222111000FFFEEEDDDCCCBBAAA9998887776665544433;
defparam prom_inst_1.INIT_RAM_0C = 256'h999888887777666655554444333322211110000FFFFEEEDDDDCCCBBBBAAA9998;
defparam prom_inst_1.INIT_RAM_0D = 256'h5555554444443333332222221111100000FFFFFFEEEEDDDDDCCCCCBBBBAAAAA9;
defparam prom_inst_1.INIT_RAM_0E = 256'hDDDDDCCCCCCCCCCCBBBBBBBBBBAAAAAAAAA99999999888888877777776666666;
defparam prom_inst_1.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEEEEEEEEEEEEEEEEEEDDDDDDDD;
defparam prom_inst_1.INIT_RAM_10 = 256'hDDDDDDDEEEEEEEEEEEEEEEEEEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_11 = 256'h6666667777777888888899999999AAAAAAAAABBBBBBBBBBCCCCCCCCCCCDDDDDD;
defparam prom_inst_1.INIT_RAM_12 = 256'hAAAAABBBBCCCCCDDDDDEEEEFFFFFF00000111112222223333334444445555556;
defparam prom_inst_1.INIT_RAM_13 = 256'h999AAABBBBCCCDDDDEEEFFFF0000111122233334444555566667777888889999;
defparam prom_inst_1.INIT_RAM_14 = 256'h344455666777888999AAABBCCCDDDEEEFFF00011122233334445556667778888;
defparam prom_inst_1.INIT_RAM_15 = 256'hAAABBCCDDDEEFF0001122233445556677788999AABBBCCDDDEEEFF0001112233;
defparam prom_inst_1.INIT_RAM_16 = 256'hCCDDEEFF001122334445566778899AABBCCDDDEEFF0011222334455666778899;
defparam prom_inst_1.INIT_RAM_17 = 256'hABBCCDDEEF0011223344556778899AABBCCDDEEFF0112233445566778899AABB;
defparam prom_inst_1.INIT_RAM_18 = 256'h55677889AABBCDDEEF00112334456677889AABBCCDEEFF001223344566778899;
defparam prom_inst_1.INIT_RAM_19 = 256'hDDEEF0012234456678899ABBCDDEFF0012234455677899AABCCDEEFF01122344;
defparam prom_inst_1.INIT_RAM_1A = 256'h123445667889AABCCDEFF011233455677899ABBCDDEFF011233455677899ABBC;
defparam prom_inst_1.INIT_RAM_1B = 256'h45667889ABBCDDEF00123345567889AABCCDEFF01123445667889ABBCDDEFF01;
defparam prom_inst_1.INIT_RAM_1C = 256'h5667899ABCCDEFF0122345567789AABCDDEF00123345667889ABBCDEEF001233;
defparam prom_inst_1.INIT_RAM_1D = 256'h45667899ABCDDEF0012334567789AABCDDEF0012334566789AABCDDEF0012334;
defparam prom_inst_1.INIT_RAM_1E = 256'h2345667899ABCDDEF0012344567789ABBCDEEF0122345567899ABCCDEFF01233;
defparam prom_inst_1.INIT_RAM_1F = 256'h012334567789AABCDEEF0122345567899ABCDDEF0012344567789ABBCDEFF012;
defparam prom_inst_1.INIT_RAM_20 = 256'hEF0012344567789ABBCDEFF0122345667899ABCDDEF0112344567889ABCCDEFF;
defparam prom_inst_1.INIT_RAM_21 = 256'hCDEFF0123345667899ABCDDEF0012344567789ABBCDEEF0122345567899ABCDD;
defparam prom_inst_1.INIT_RAM_22 = 256'hCCDEFF0122345567889ABBCDEFF0122345567889ABBCDEFF0122345567899ABC;
defparam prom_inst_1.INIT_RAM_23 = 256'hCDEEF01123445667899ABCCDEFF0122344567789AABCDDEF00123345667899AB;
defparam prom_inst_1.INIT_RAM_24 = 256'hF001223445667899ABBCDEEF00122345567789AABCCDEFF01123445667899ABC;
defparam prom_inst_1.INIT_RAM_25 = 256'h445667889AABCCDEEF001223445667889AABCCDEEF001223455677899ABBCDDE;
defparam prom_inst_1.INIT_RAM_26 = 256'hBCDDEEF00112334556678899ABBCDDEFF0012234455677899ABBCDDEEF001223;
defparam prom_inst_1.INIT_RAM_27 = 256'h6778899ABBCCDDEEF001122344556778899ABBCCDEEFF00122334556678899AB;
defparam prom_inst_1.INIT_RAM_28 = 256'h45566778899AABBCCDDEEFF0012233445566778899ABBCCDDEEFF01122334455;
defparam prom_inst_1.INIT_RAM_29 = 256'h67788899AABBCCCDDEEFF0011122334455667788999AABBCCDDEEFF001122334;
defparam prom_inst_1.INIT_RAM_2A = 256'hCDDDEEFFF0001122233444556667788899AAABBCCCDDEEFFF001112233445556;
defparam prom_inst_1.INIT_RAM_2B = 256'h777888999AAABBBBCCCDDDEEEFFF00011122233344455566777888999AABBBCC;
defparam prom_inst_1.INIT_RAM_2C = 256'h6666777788889999AAAABBBBCCCCDDDDEEEFFFF0000111222233344445556667;
defparam prom_inst_1.INIT_RAM_2D = 256'hAAAAAAABBBBBBCCCCCCDDDDDEEEEEEFFFFF00000111112222233334444455556;
defparam prom_inst_1.INIT_RAM_2E = 256'h2222223333333333344444444455555555566666666777777778888888999999;
defparam prom_inst_1.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000111111111111111112222222;
defparam prom_inst_1.INIT_RAM_30 = 256'h2222221111111111111111100000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_31 = 256'h9999988888887777777766666666555555555444444444333333333332222222;
defparam prom_inst_1.INIT_RAM_32 = 256'h5555444443333222221111100000FFFFFEEEEEEDDDDDCCCCCCBBBBBBAAAAAAA9;
defparam prom_inst_1.INIT_RAM_33 = 256'h666555444433322221110000FFFFEEEDDDDCCCCBBBBAAAA99998888777766666;
defparam prom_inst_1.INIT_RAM_34 = 256'hCBBBAA99988877766555444333222111000FFFEEEDDDCCCBBBBAAA9998887777;
defparam prom_inst_1.INIT_RAM_35 = 256'h55544332211100FFFEEDDCCCBBAAA9988877666554443322211000FFFEEDDDCC;
defparam prom_inst_1.INIT_RAM_36 = 256'h33221100FFEEDDCCBBAA9998877665544332211100FFEEDDCCCBBAA998887766;
defparam prom_inst_1.INIT_RAM_37 = 256'h5443322110FFEEDDCCBBA9988776655443322100FFEEDDCCBBAA998877665544;
defparam prom_inst_1.INIT_RAM_38 = 256'hA99887665543322100FFEEDCCBBA998877655443221100FEEDDCCBBA99887765;
defparam prom_inst_1.INIT_RAM_39 = 256'h22100FEEDDCBBA9987765544322100FFEDDCBBA99887665543321100FEEDDCBB;
defparam prom_inst_1.INIT_RAM_3A = 256'hDDCBBA998776554322100FEEDCCBAA988766544322100FEEDCCBAA9887665443;
defparam prom_inst_1.INIT_RAM_3B = 256'hBA99876654432110FFEDCCBAA98776554322100FEEDCBBA998766544322100FE;
defparam prom_inst_1.INIT_RAM_3C = 256'hA99876654332100FEDDCBAA9877654432210FFEDCCBA99876654432110FEEDCC;
defparam prom_inst_1.INIT_RAM_3D = 256'hBA9987655432210FFEDCBBA9887655432210FFEDCBBA9887655432210FFEDCCB;
defparam prom_inst_1.INIT_RAM_3E = 256'hDCBA9987655432210FEEDCBBA9877654432100FEDDCBA9987665433210FFEDCC;
defparam prom_inst_1.INIT_RAM_3F = 256'hFEDCCBA9887654432110FEDDCBA9987665432210FFEDCBBA9877654432100FED;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[27:0],dout[11:8]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 4;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'h332222222222222222222221111111111111111111100000000000000000000F;
defparam prom_inst_2.INIT_RAM_01 = 256'h6666555555555555555555555444444444444444444444333333333333333333;
defparam prom_inst_2.INIT_RAM_02 = 256'h9999998888888888888888888887777777777777777777776666666666666666;
defparam prom_inst_2.INIT_RAM_03 = 256'hCCCCCBBBBBBBBBBBBBBBBBBBBBBAAAAAAAAAAAAAAAAAAAAA9999999999999999;
defparam prom_inst_2.INIT_RAM_04 = 256'hFEEEEEEEEEEEEEEEEEEEEEEEDDDDDDDDDDDDDDDDDDDDDDDCCCCCCCCCCCCCCCCC;
defparam prom_inst_2.INIT_RAM_05 = 256'h111111111111111111000000000000000000000000FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_06 = 256'h4444444333333333333333333333333332222222222222222222222222111111;
defparam prom_inst_2.INIT_RAM_07 = 256'h6666666666666666655555555555555555555555555554444444444444444444;
defparam prom_inst_2.INIT_RAM_08 = 256'h8888888888888888888888777777777777777777777777777777766666666666;
defparam prom_inst_2.INIT_RAM_09 = 256'hAAAAAAAAAAAAAAAAAAAAA9999999999999999999999999999999999888888888;
defparam prom_inst_2.INIT_RAM_0A = 256'hCCCCCCCCCBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBAAAAAAAAAAAAAAA;
defparam prom_inst_2.INIT_RAM_0B = 256'hDDDDDDDDDDDDDDDDDDDDDDDDDDDDCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCC;
defparam prom_inst_2.INIT_RAM_0C = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEDDDDDDDDDDDDDDDDDDDDDDDDD;
defparam prom_inst_2.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam prom_inst_2.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_12 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_13 = 256'hDDDDDDDDDDDDDDDDDDDDDDDDEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam prom_inst_2.INIT_RAM_14 = 256'hCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCDDDDDDDDDDDDDDDDDDDDDDDDDDDDD;
defparam prom_inst_2.INIT_RAM_15 = 256'hAAAAAAAAAAAAAABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBCCCCCCCCCC;
defparam prom_inst_2.INIT_RAM_16 = 256'h888888889999999999999999999999999999999999AAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_2.INIT_RAM_17 = 256'h6666666666777777777777777777777777777777788888888888888888888888;
defparam prom_inst_2.INIT_RAM_18 = 256'h4444444444444444445555555555555555555555555555666666666666666666;
defparam prom_inst_2.INIT_RAM_19 = 256'h1111122222222222222222222222223333333333333333333333333344444444;
defparam prom_inst_2.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFF0000000000000000000000001111111111111111111;
defparam prom_inst_2.INIT_RAM_1B = 256'hCCCCCCCCCCCCCCCCDDDDDDDDDDDDDDDDDDDDDDDEEEEEEEEEEEEEEEEEEEEEEEFF;
defparam prom_inst_2.INIT_RAM_1C = 256'h999999999999999AAAAAAAAAAAAAAAAAAAAABBBBBBBBBBBBBBBBBBBBBBCCCCCC;
defparam prom_inst_2.INIT_RAM_1D = 256'h6666666666666667777777777777777777778888888888888888888889999999;
defparam prom_inst_2.INIT_RAM_1E = 256'h3333333333333333344444444444444444444455555555555555555555566666;
defparam prom_inst_2.INIT_RAM_1F = 256'h0000000000000000000011111111111111111111222222222222222222222333;
defparam prom_inst_2.INIT_RAM_20 = 256'hCCDDDDDDDDDDDDDDDDDDDDDEEEEEEEEEEEEEEEEEEEEFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_21 = 256'h99999AAAAAAAAAAAAAAAAAAAABBBBBBBBBBBBBBBBBBBBBCCCCCCCCCCCCCCCCCC;
defparam prom_inst_2.INIT_RAM_22 = 256'h6666667777777777777777777778888888888888888888889999999999999999;
defparam prom_inst_2.INIT_RAM_23 = 256'h3333344444444444444444444445555555555555555555556666666666666666;
defparam prom_inst_2.INIT_RAM_24 = 256'h0111111111111111111111112222222222222222222222233333333333333333;
defparam prom_inst_2.INIT_RAM_25 = 256'hEEEEEEEEEEEEEEEEEEFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000;
defparam prom_inst_2.INIT_RAM_26 = 256'hBBBBBBBCCCCCCCCCCCCCCCCCCCCCCCCCCDDDDDDDDDDDDDDDDDDDDDDDDDEEEEEE;
defparam prom_inst_2.INIT_RAM_27 = 256'h99999999999999999AAAAAAAAAAAAAAAAAAAAAAAAAAAABBBBBBBBBBBBBBBBBBB;
defparam prom_inst_2.INIT_RAM_28 = 256'h7777777777777777777777788888888888888888888888888888899999999999;
defparam prom_inst_2.INIT_RAM_29 = 256'h5555555555555555555556666666666666666666666666666666666777777777;
defparam prom_inst_2.INIT_RAM_2A = 256'h3333333334444444444444444444444444444444444444444555555555555555;
defparam prom_inst_2.INIT_RAM_2B = 256'h2222222222222222222222222222333333333333333333333333333333333333;
defparam prom_inst_2.INIT_RAM_2C = 256'h1111111111111111111111111111111111111112222222222222222222222222;
defparam prom_inst_2.INIT_RAM_2D = 256'h0000000000000000000000000000000000011111111111111111111111111111;
defparam prom_inst_2.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_32 = 256'h1111111111111111111111111111000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_33 = 256'h2222222222222222222222221111111111111111111111111111111111111111;
defparam prom_inst_2.INIT_RAM_34 = 256'h3333333333333333333333333333333333322222222222222222222222222222;
defparam prom_inst_2.INIT_RAM_35 = 256'h5555555555555544444444444444444444444444444444444444443333333333;
defparam prom_inst_2.INIT_RAM_36 = 256'h7777777766666666666666666666666666666666665555555555555555555555;
defparam prom_inst_2.INIT_RAM_37 = 256'h9999999999888888888888888888888888888888777777777777777777777777;
defparam prom_inst_2.INIT_RAM_38 = 256'hBBBBBBBBBBBBBBBBBBAAAAAAAAAAAAAAAAAAAAAAAAAAAA999999999999999999;
defparam prom_inst_2.INIT_RAM_39 = 256'hEEEEEDDDDDDDDDDDDDDDDDDDDDDDDDCCCCCCCCCCCCCCCCCCCCCCCCCCBBBBBBBB;
defparam prom_inst_2.INIT_RAM_3A = 256'h000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFEEEEEEEEEEEEEEEEEEE;
defparam prom_inst_2.INIT_RAM_3B = 256'h3333333333333333222222222222222222222221111111111111111111111100;
defparam prom_inst_2.INIT_RAM_3C = 256'h6666666666666665555555555555555555554444444444444444444444333333;
defparam prom_inst_2.INIT_RAM_3D = 256'h9999999999999998888888888888888888887777777777777777777776666666;
defparam prom_inst_2.INIT_RAM_3E = 256'hCCCCCCCCCCCCCCCCCBBBBBBBBBBBBBBBBBBBBBAAAAAAAAAAAAAAAAAAAA999999;
defparam prom_inst_2.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFEEEEEEEEEEEEEEEEEEEEDDDDDDDDDDDDDDDDDDDDDCCC;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[29:0],dout[13:12]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({gw_gnd,ad[11:0],gw_gnd})
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 2;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9;
defparam prom_inst_3.INIT_RAM_01 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_3.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_3.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_0D = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAABFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_0E = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_3.INIT_RAM_0F = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_3.INIT_RAM_10 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
defparam prom_inst_3.INIT_RAM_11 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
defparam prom_inst_3.INIT_RAM_12 = 256'h0000000000000000000005555555555555555555555555555555555555555555;
defparam prom_inst_3.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_1D = 256'h5555555555555555555555555555555555555555554000000000000000000000;
defparam prom_inst_3.INIT_RAM_1E = 256'h5555555555555555555555555555555555555555555555555555555555555555;
defparam prom_inst_3.INIT_RAM_1F = 256'h5555555555555555555555555555555555555555555555555555555555555555;

endmodule //rom_sine
