`timescale 1ns/1ps

module dac_engine_tb();
    
    reg clk;
    reg rst_n;
    reg enable;
    reg [31:0] freq;
    reg [15:0] phase_offset;
    reg [15:0] amplitude;
    reg wr_en;
    reg [8:0] wr_addr;
    reg [15:0] wr_data;
    reg high_quality_mode;
    
    wire [15:0] dac_out;
    
    integer i, output_file;
    
    dac_engine u_dds (
        .clk(clk),
        .rst_n(rst_n),
        .dds_enable(enable),
        .frequency(freq),
        .amplitude(amplitude),
        .phase_offset(phase_offset),
        .wave_wr_en(wr_en),
        .wave_addr(wr_addr),
        .wave_data(wr_data),
        .high_quality_mode(high_quality_mode),
        .dac_out(dac_out)
    );
    
    // Clock generation
    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end
    
    initial begin
        // Initialize
        rst_n = 0;
        enable = 0;
        freq = 0;
        phase_offset = 0;
        amplitude = 16'h7FFF;
        high_quality_mode = 0;
        wr_en = 0;
        wr_addr = 0;
        wr_data = 0;
        
        #100;
        rst_n = 1;
        #100;
        
        $display("=== Final DDS Verification Test ===");
        
        // 1. Initialize complete sine wave
        $display("1. Initializing 512-point sine wave...");
        for (i = 0; i < 512; i = i + 1) begin
            @(posedge clk);
            wr_en = 1;
            wr_addr = i;
            wr_data = $rtoi(32767.0 * $sin(2.0 * 3.1415926 * i / 512.0));
        end
        @(posedge clk);
        wr_en = 0;
        #100;
        
        // 2. Test normal mode (linear interpolation)
        $display("2. Testing normal mode (linear interpolation)...");
        freq = 32'h20000000; // Medium frequency
        enable = 1;
        high_quality_mode = 0;
        
        output_file = $fopen("normal_mode_output.txt", "w");
        for (i = 0; i < 100; i = i + 1) begin
            @(posedge clk);
            $fwrite(output_file, "%d\n", $signed(dac_out));
        end
        $fclose(output_file);
        enable = 0;
        #100;
        
        // 3. Test high quality mode (cubic interpolation)
        $display("3. Testing high quality mode (cubic interpolation)...");
        freq = 32'h20000000;
        enable = 1;
        high_quality_mode = 1;
        
        output_file = $fopen("high_quality_output.txt", "w");
        for (i = 0; i < 100; i = i + 1) begin
            @(posedge clk);
            $fwrite(output_file, "%d\n", $signed(dac_out));
        end
        $fclose(output_file);
        enable = 0;
        #100;
        
        // 4. Test frequency response
        $display("4. Testing frequency response...");
        enable = 1;
        high_quality_mode = 1;
        
        // Sweep frequencies
        freq = 32'h08000000; // Low frequency
        #1000;
        
        freq = 32'h20000000; // Medium frequency  
        #1000;
        
        freq = 32'h40000000; // High frequency
        #1000;
        
        enable = 0;
        #100;
        
        $display("=== All Verification Tests Completed Successfully ===");
        $display("DDS System is fully functional!");
        $finish;
    end
    
    // Monitor for real-time verification
    always @(posedge clk) begin
        if (enable && $time > 1000) begin
            // Check for valid output range
            if ($signed(dac_out) > 32767 || $signed(dac_out) < -32768) begin
                $display("WARNING: Output out of range: %d", $signed(dac_out));
            end
        end
    end
    
    initial begin
        $dumpfile("dac_engine_tb.vcd");
        $dumpvars(0, dac_engine_tb);
    end

endmodule