module triangular_rom_a8d8(
	addr,
	clk, 
	q
);	

	parameter DATA_WIDTH=8;
	parameter ADDR_WIDTH=8;

	input clk;
	input [(ADDR_WIDTH-1):0] addr;
	output reg [(DATA_WIDTH-1):0] q;
	


	// Declare the ROM variable
	reg [DATA_WIDTH-1:0] rom[2**ADDR_WIDTH-1:0];

	initial begin
		rom[000] = 8'h0; 
		rom[001] = 8'h2; 
		rom[002] = 8'h4; 
		rom[003] = 8'h6; 
		rom[004] = 8'h8; 
		rom[005] = 8'ha; 
		rom[006] = 8'hc; 
		rom[007] = 8'he; 
		rom[008] = 8'h10; 
		rom[009] = 8'h12; 
		rom[010] = 8'h14; 
		rom[011] = 8'h16; 
		rom[012] = 8'h18; 
		rom[013] = 8'h1a; 
		rom[014] = 8'h1c; 
		rom[015] = 8'h1e; 
		rom[016] = 8'h20; 
		rom[017] = 8'h22; 
		rom[018] = 8'h24; 
		rom[019] = 8'h26; 
		rom[020] = 8'h28; 
		rom[021] = 8'h2a; 
		rom[022] = 8'h2c; 
		rom[023] = 8'h2e; 
		rom[024] = 8'h30; 
		rom[025] = 8'h32; 
		rom[026] = 8'h34; 
		rom[027] = 8'h36; 
		rom[028] = 8'h38; 
		rom[029] = 8'h3a; 
		rom[030] = 8'h3c; 
		rom[031] = 8'h3e; 
		rom[032] = 8'h40; 
		rom[033] = 8'h42; 
		rom[034] = 8'h44; 
		rom[035] = 8'h46; 
		rom[036] = 8'h48; 
		rom[037] = 8'h4a; 
		rom[038] = 8'h4c; 
		rom[039] = 8'h4e; 
		rom[040] = 8'h50; 
		rom[041] = 8'h52; 
		rom[042] = 8'h54; 
		rom[043] = 8'h56; 
		rom[044] = 8'h58; 
		rom[045] = 8'h5a; 
		rom[046] = 8'h5c; 
		rom[047] = 8'h5e; 
		rom[048] = 8'h60; 
		rom[049] = 8'h62; 
		rom[050] = 8'h64; 
		rom[051] = 8'h66; 
		rom[052] = 8'h68; 
		rom[053] = 8'h6a; 
		rom[054] = 8'h6c; 
		rom[055] = 8'h6e; 
		rom[056] = 8'h70; 
		rom[057] = 8'h72; 
		rom[058] = 8'h74; 
		rom[059] = 8'h76; 
		rom[060] = 8'h78; 
		rom[061] = 8'h7a; 
		rom[062] = 8'h7c; 
		rom[063] = 8'h7e; 
		rom[064] = 8'h80; 
		rom[065] = 8'h81; 
		rom[066] = 8'h83; 
		rom[067] = 8'h85; 
		rom[068] = 8'h87; 
		rom[069] = 8'h89; 
		rom[070] = 8'h8b; 
		rom[071] = 8'h8d; 
		rom[072] = 8'h8f; 
		rom[073] = 8'h91; 
		rom[074] = 8'h93; 
		rom[075] = 8'h95; 
		rom[076] = 8'h97; 
		rom[077] = 8'h99; 
		rom[078] = 8'h9b; 
		rom[079] = 8'h9d; 
		rom[080] = 8'h9f; 
		rom[081] = 8'ha1; 
		rom[082] = 8'ha3; 
		rom[083] = 8'ha5; 
		rom[084] = 8'ha7; 
		rom[085] = 8'ha9; 
		rom[086] = 8'hab; 
		rom[087] = 8'had; 
		rom[088] = 8'haf; 
		rom[089] = 8'hb1; 
		rom[090] = 8'hb3; 
		rom[091] = 8'hb5; 
		rom[092] = 8'hb7; 
		rom[093] = 8'hb9; 
		rom[094] = 8'hbb; 
		rom[095] = 8'hbd; 
		rom[096] = 8'hbf; 
		rom[097] = 8'hc1; 
		rom[098] = 8'hc3; 
		rom[099] = 8'hc5; 
		rom[100] = 8'hc7; 
		rom[101] = 8'hc9; 
		rom[102] = 8'hcb; 
		rom[103] = 8'hcd; 
		rom[104] = 8'hcf; 
		rom[105] = 8'hd1; 
		rom[106] = 8'hd3; 
		rom[107] = 8'hd5; 
		rom[108] = 8'hd7; 
		rom[109] = 8'hd9; 
		rom[110] = 8'hdb; 
		rom[111] = 8'hdd; 
		rom[112] = 8'hdf; 
		rom[113] = 8'he1; 
		rom[114] = 8'he3; 
		rom[115] = 8'he5; 
		rom[116] = 8'he7; 
		rom[117] = 8'he9; 
		rom[118] = 8'heb; 
		rom[119] = 8'hed; 
		rom[120] = 8'hef; 
		rom[121] = 8'hf1; 
		rom[122] = 8'hf3; 
		rom[123] = 8'hf5; 
		rom[124] = 8'hf7; 
		rom[125] = 8'hf9; 
		rom[126] = 8'hfb; 
		rom[127] = 8'hfd; 
		rom[128] = 8'hff; 
		rom[129] = 8'hfd; 
		rom[130] = 8'hfb; 
		rom[131] = 8'hf9; 
		rom[132] = 8'hf7; 
		rom[133] = 8'hf5; 
		rom[134] = 8'hf3; 
		rom[135] = 8'hf1; 
		rom[136] = 8'hef; 
		rom[137] = 8'hed; 
		rom[138] = 8'heb; 
		rom[139] = 8'he9; 
		rom[140] = 8'he7; 
		rom[141] = 8'he5; 
		rom[142] = 8'he3; 
		rom[143] = 8'he1; 
		rom[144] = 8'hdf; 
		rom[145] = 8'hdd; 
		rom[146] = 8'hdb; 
		rom[147] = 8'hd9; 
		rom[148] = 8'hd7; 
		rom[149] = 8'hd5; 
		rom[150] = 8'hd3; 
		rom[151] = 8'hd1; 
		rom[152] = 8'hcf; 
		rom[153] = 8'hcd; 
		rom[154] = 8'hcb; 
		rom[155] = 8'hc9; 
		rom[156] = 8'hc7; 
		rom[157] = 8'hc5; 
		rom[158] = 8'hc3; 
		rom[159] = 8'hc1; 
		rom[160] = 8'hbf; 
		rom[161] = 8'hbd; 
		rom[162] = 8'hbb; 
		rom[163] = 8'hb9; 
		rom[164] = 8'hb7; 
		rom[165] = 8'hb5; 
		rom[166] = 8'hb3; 
		rom[167] = 8'hb1; 
		rom[168] = 8'haf; 
		rom[169] = 8'had; 
		rom[170] = 8'hab; 
		rom[171] = 8'ha9; 
		rom[172] = 8'ha7; 
		rom[173] = 8'ha5; 
		rom[174] = 8'ha3; 
		rom[175] = 8'ha1; 
		rom[176] = 8'h9f; 
		rom[177] = 8'h9d; 
		rom[178] = 8'h9b; 
		rom[179] = 8'h99; 
		rom[180] = 8'h97; 
		rom[181] = 8'h95; 
		rom[182] = 8'h93; 
		rom[183] = 8'h91; 
		rom[184] = 8'h8f; 
		rom[185] = 8'h8d; 
		rom[186] = 8'h8b; 
		rom[187] = 8'h89; 
		rom[188] = 8'h87; 
		rom[189] = 8'h85; 
		rom[190] = 8'h83; 
		rom[191] = 8'h81; 
		rom[192] = 8'h80; 
		rom[193] = 8'h7e; 
		rom[194] = 8'h7c; 
		rom[195] = 8'h7a; 
		rom[196] = 8'h78; 
		rom[197] = 8'h76; 
		rom[198] = 8'h74; 
		rom[199] = 8'h72; 
		rom[200] = 8'h70; 
		rom[201] = 8'h6e; 
		rom[202] = 8'h6c; 
		rom[203] = 8'h6a; 
		rom[204] = 8'h68; 
		rom[205] = 8'h66; 
		rom[206] = 8'h64; 
		rom[207] = 8'h62; 
		rom[208] = 8'h60; 
		rom[209] = 8'h5e; 
		rom[210] = 8'h5c; 
		rom[211] = 8'h5a; 
		rom[212] = 8'h58; 
		rom[213] = 8'h56; 
		rom[214] = 8'h54; 
		rom[215] = 8'h52; 
		rom[216] = 8'h50; 
		rom[217] = 8'h4e; 
		rom[218] = 8'h4c; 
		rom[219] = 8'h4a; 
		rom[220] = 8'h48; 
		rom[221] = 8'h46; 
		rom[222] = 8'h44; 
		rom[223] = 8'h42; 
		rom[224] = 8'h40; 
		rom[225] = 8'h3e; 
		rom[226] = 8'h3c; 
		rom[227] = 8'h3a; 
		rom[228] = 8'h38; 
		rom[229] = 8'h36; 
		rom[230] = 8'h34; 
		rom[231] = 8'h32; 
		rom[232] = 8'h30; 
		rom[233] = 8'h2e; 
		rom[234] = 8'h2c; 
		rom[235] = 8'h2a; 
		rom[236] = 8'h28; 
		rom[237] = 8'h26; 
		rom[238] = 8'h24; 
		rom[239] = 8'h22; 
		rom[240] = 8'h20; 
		rom[241] = 8'h1e; 
		rom[242] = 8'h1c; 
		rom[243] = 8'h1a; 
		rom[244] = 8'h18; 
		rom[245] = 8'h16; 
		rom[246] = 8'h14; 
		rom[247] = 8'h12; 
		rom[248] = 8'h10; 
		rom[249] = 8'he; 
		rom[250] = 8'hc; 
		rom[251] = 8'ha; 
		rom[252] = 8'h8; 
		rom[253] = 8'h6; 
		rom[254] = 8'h4; 
		rom[255] = 8'h2; 
	end

	always @ (posedge clk)
	begin
		q <= rom[addr];
	end

endmodule
