module square_wave_rom_a8d8(
	addr,
	clk, 
	q
);	

	parameter DATA_WIDTH=8;
	parameter ADDR_WIDTH=8;

	input clk;
	input [(ADDR_WIDTH-1):0] addr;
	output reg [(DATA_WIDTH-1):0] q;
	


	// Declare the ROM variable
	reg [DATA_WIDTH-1:0] rom[2**ADDR_WIDTH-1:0];

	initial begin
		rom[000] = 8'hff; 
		rom[001] = 8'hff; 
		rom[002] = 8'hff; 
		rom[003] = 8'hff; 
		rom[004] = 8'hff; 
		rom[005] = 8'hff; 
		rom[006] = 8'hff; 
		rom[007] = 8'hff; 
		rom[008] = 8'hff; 
		rom[009] = 8'hff; 
		rom[010] = 8'hff; 
		rom[011] = 8'hff; 
		rom[012] = 8'hff; 
		rom[013] = 8'hff; 
		rom[014] = 8'hff; 
		rom[015] = 8'hff; 
		rom[016] = 8'hff; 
		rom[017] = 8'hff; 
		rom[018] = 8'hff; 
		rom[019] = 8'hff; 
		rom[020] = 8'hff; 
		rom[021] = 8'hff; 
		rom[022] = 8'hff; 
		rom[023] = 8'hff; 
		rom[024] = 8'hff; 
		rom[025] = 8'hff; 
		rom[026] = 8'hff; 
		rom[027] = 8'hff; 
		rom[028] = 8'hff; 
		rom[029] = 8'hff; 
		rom[030] = 8'hff; 
		rom[031] = 8'hff; 
		rom[032] = 8'hff; 
		rom[033] = 8'hff; 
		rom[034] = 8'hff; 
		rom[035] = 8'hff; 
		rom[036] = 8'hff; 
		rom[037] = 8'hff; 
		rom[038] = 8'hff; 
		rom[039] = 8'hff; 
		rom[040] = 8'hff; 
		rom[041] = 8'hff; 
		rom[042] = 8'hff; 
		rom[043] = 8'hff; 
		rom[044] = 8'hff; 
		rom[045] = 8'hff; 
		rom[046] = 8'hff; 
		rom[047] = 8'hff; 
		rom[048] = 8'hff; 
		rom[049] = 8'hff; 
		rom[050] = 8'hff; 
		rom[051] = 8'hff; 
		rom[052] = 8'hff; 
		rom[053] = 8'hff; 
		rom[054] = 8'hff; 
		rom[055] = 8'hff; 
		rom[056] = 8'hff; 
		rom[057] = 8'hff; 
		rom[058] = 8'hff; 
		rom[059] = 8'hff; 
		rom[060] = 8'hff; 
		rom[061] = 8'hff; 
		rom[062] = 8'hff; 
		rom[063] = 8'hff; 
		rom[064] = 8'hff; 
		rom[065] = 8'hff; 
		rom[066] = 8'hff; 
		rom[067] = 8'hff; 
		rom[068] = 8'hff; 
		rom[069] = 8'hff; 
		rom[070] = 8'hff; 
		rom[071] = 8'hff; 
		rom[072] = 8'hff; 
		rom[073] = 8'hff; 
		rom[074] = 8'hff; 
		rom[075] = 8'hff; 
		rom[076] = 8'hff; 
		rom[077] = 8'hff; 
		rom[078] = 8'hff; 
		rom[079] = 8'hff; 
		rom[080] = 8'hff; 
		rom[081] = 8'hff; 
		rom[082] = 8'hff; 
		rom[083] = 8'hff; 
		rom[084] = 8'hff; 
		rom[085] = 8'hff; 
		rom[086] = 8'hff; 
		rom[087] = 8'hff; 
		rom[088] = 8'hff; 
		rom[089] = 8'hff; 
		rom[090] = 8'hff; 
		rom[091] = 8'hff; 
		rom[092] = 8'hff; 
		rom[093] = 8'hff; 
		rom[094] = 8'hff; 
		rom[095] = 8'hff; 
		rom[096] = 8'hff; 
		rom[097] = 8'hff; 
		rom[098] = 8'hff; 
		rom[099] = 8'hff; 
		rom[100] = 8'hff; 
		rom[101] = 8'hff; 
		rom[102] = 8'hff; 
		rom[103] = 8'hff; 
		rom[104] = 8'hff; 
		rom[105] = 8'hff; 
		rom[106] = 8'hff; 
		rom[107] = 8'hff; 
		rom[108] = 8'hff; 
		rom[109] = 8'hff; 
		rom[110] = 8'hff; 
		rom[111] = 8'hff; 
		rom[112] = 8'hff; 
		rom[113] = 8'hff; 
		rom[114] = 8'hff; 
		rom[115] = 8'hff; 
		rom[116] = 8'hff; 
		rom[117] = 8'hff; 
		rom[118] = 8'hff; 
		rom[119] = 8'hff; 
		rom[120] = 8'hff; 
		rom[121] = 8'hff; 
		rom[122] = 8'hff; 
		rom[123] = 8'hff; 
		rom[124] = 8'hff; 
		rom[125] = 8'hff; 
		rom[126] = 8'hff; 
		rom[127] = 8'hff; 
		rom[128] = 8'h0; 
		rom[129] = 8'h0; 
		rom[130] = 8'h0; 
		rom[131] = 8'h0; 
		rom[132] = 8'h0; 
		rom[133] = 8'h0; 
		rom[134] = 8'h0; 
		rom[135] = 8'h0; 
		rom[136] = 8'h0; 
		rom[137] = 8'h0; 
		rom[138] = 8'h0; 
		rom[139] = 8'h0; 
		rom[140] = 8'h0; 
		rom[141] = 8'h0; 
		rom[142] = 8'h0; 
		rom[143] = 8'h0; 
		rom[144] = 8'h0; 
		rom[145] = 8'h0; 
		rom[146] = 8'h0; 
		rom[147] = 8'h0; 
		rom[148] = 8'h0; 
		rom[149] = 8'h0; 
		rom[150] = 8'h0; 
		rom[151] = 8'h0; 
		rom[152] = 8'h0; 
		rom[153] = 8'h0; 
		rom[154] = 8'h0; 
		rom[155] = 8'h0; 
		rom[156] = 8'h0; 
		rom[157] = 8'h0; 
		rom[158] = 8'h0; 
		rom[159] = 8'h0; 
		rom[160] = 8'h0; 
		rom[161] = 8'h0; 
		rom[162] = 8'h0; 
		rom[163] = 8'h0; 
		rom[164] = 8'h0; 
		rom[165] = 8'h0; 
		rom[166] = 8'h0; 
		rom[167] = 8'h0; 
		rom[168] = 8'h0; 
		rom[169] = 8'h0; 
		rom[170] = 8'h0; 
		rom[171] = 8'h0; 
		rom[172] = 8'h0; 
		rom[173] = 8'h0; 
		rom[174] = 8'h0; 
		rom[175] = 8'h0; 
		rom[176] = 8'h0; 
		rom[177] = 8'h0; 
		rom[178] = 8'h0; 
		rom[179] = 8'h0; 
		rom[180] = 8'h0; 
		rom[181] = 8'h0; 
		rom[182] = 8'h0; 
		rom[183] = 8'h0; 
		rom[184] = 8'h0; 
		rom[185] = 8'h0; 
		rom[186] = 8'h0; 
		rom[187] = 8'h0; 
		rom[188] = 8'h0; 
		rom[189] = 8'h0; 
		rom[190] = 8'h0; 
		rom[191] = 8'h0; 
		rom[192] = 8'h0; 
		rom[193] = 8'h0; 
		rom[194] = 8'h0; 
		rom[195] = 8'h0; 
		rom[196] = 8'h0; 
		rom[197] = 8'h0; 
		rom[198] = 8'h0; 
		rom[199] = 8'h0; 
		rom[200] = 8'h0; 
		rom[201] = 8'h0; 
		rom[202] = 8'h0; 
		rom[203] = 8'h0; 
		rom[204] = 8'h0; 
		rom[205] = 8'h0; 
		rom[206] = 8'h0; 
		rom[207] = 8'h0; 
		rom[208] = 8'h0; 
		rom[209] = 8'h0; 
		rom[210] = 8'h0; 
		rom[211] = 8'h0; 
		rom[212] = 8'h0; 
		rom[213] = 8'h0; 
		rom[214] = 8'h0; 
		rom[215] = 8'h0; 
		rom[216] = 8'h0; 
		rom[217] = 8'h0; 
		rom[218] = 8'h0; 
		rom[219] = 8'h0; 
		rom[220] = 8'h0; 
		rom[221] = 8'h0; 
		rom[222] = 8'h0; 
		rom[223] = 8'h0; 
		rom[224] = 8'h0; 
		rom[225] = 8'h0; 
		rom[226] = 8'h0; 
		rom[227] = 8'h0; 
		rom[228] = 8'h0; 
		rom[229] = 8'h0; 
		rom[230] = 8'h0; 
		rom[231] = 8'h0; 
		rom[232] = 8'h0; 
		rom[233] = 8'h0; 
		rom[234] = 8'h0; 
		rom[235] = 8'h0; 
		rom[236] = 8'h0; 
		rom[237] = 8'h0; 
		rom[238] = 8'h0; 
		rom[239] = 8'h0; 
		rom[240] = 8'h0; 
		rom[241] = 8'h0; 
		rom[242] = 8'h0; 
		rom[243] = 8'h0; 
		rom[244] = 8'h0; 
		rom[245] = 8'h0; 
		rom[246] = 8'h0; 
		rom[247] = 8'h0; 
		rom[248] = 8'h0; 
		rom[249] = 8'h0; 
		rom[250] = 8'h0; 
		rom[251] = 8'h0; 
		rom[252] = 8'h0; 
		rom[253] = 8'h0; 
		rom[254] = 8'h0; 
		rom[255] = 8'h0; 
	end

	always @ (posedge clk)
	begin
		q <= rom[addr];
	end

endmodule
