// -----------------------------------------------------
// 8-bit x 256 sawtooth ROM (0x00 .. 0xFF), table-assigned
// Interface identical to sin_rom_a8d8
// -----------------------------------------------------
module saw_rom_a8d8(
    addr,
    clk, 
    q
);  

    parameter DATA_WIDTH=8;
    parameter ADDR_WIDTH=8;

    input clk;
    input [(ADDR_WIDTH-1):0] addr;
    output reg [(DATA_WIDTH-1):0] q;

    // Declare the ROM variable
    reg [DATA_WIDTH-1:0] rom[2**ADDR_WIDTH-1:0];

    initial begin
        rom[000] = 8'h00; 
        rom[001] = 8'h01; 
        rom[002] = 8'h02; 
        rom[003] = 8'h03; 
        rom[004] = 8'h04; 
        rom[005] = 8'h05; 
        rom[006] = 8'h06; 
        rom[007] = 8'h07; 
        rom[008] = 8'h08; 
        rom[009] = 8'h09; 
        rom[010] = 8'h0a; 
        rom[011] = 8'h0b; 
        rom[012] = 8'h0c; 
        rom[013] = 8'h0d; 
        rom[014] = 8'h0e; 
        rom[015] = 8'h0f; 
        rom[016] = 8'h10; 
        rom[017] = 8'h11; 
        rom[018] = 8'h12; 
        rom[019] = 8'h13; 
        rom[020] = 8'h14; 
        rom[021] = 8'h15; 
        rom[022] = 8'h16; 
        rom[023] = 8'h17; 
        rom[024] = 8'h18; 
        rom[025] = 8'h19; 
        rom[026] = 8'h1a; 
        rom[027] = 8'h1b; 
        rom[028] = 8'h1c; 
        rom[029] = 8'h1d; 
        rom[030] = 8'h1e; 
        rom[031] = 8'h1f; 
        rom[032] = 8'h20; 
        rom[033] = 8'h21; 
        rom[034] = 8'h22; 
        rom[035] = 8'h23; 
        rom[036] = 8'h24; 
        rom[037] = 8'h25; 
        rom[038] = 8'h26; 
        rom[039] = 8'h27; 
        rom[040] = 8'h28; 
        rom[041] = 8'h29; 
        rom[042] = 8'h2a; 
        rom[043] = 8'h2b; 
        rom[044] = 8'h2c; 
        rom[045] = 8'h2d; 
        rom[046] = 8'h2e; 
        rom[047] = 8'h2f; 
        rom[048] = 8'h30; 
        rom[049] = 8'h31; 
        rom[050] = 8'h32; 
        rom[051] = 8'h33; 
        rom[052] = 8'h34; 
        rom[053] = 8'h35; 
        rom[054] = 8'h36; 
        rom[055] = 8'h37; 
        rom[056] = 8'h38; 
        rom[057] = 8'h39; 
        rom[058] = 8'h3a; 
        rom[059] = 8'h3b; 
        rom[060] = 8'h3c; 
        rom[061] = 8'h3d; 
        rom[062] = 8'h3e; 
        rom[063] = 8'h3f; 
        rom[064] = 8'h40; 
        rom[065] = 8'h41; 
        rom[066] = 8'h42; 
        rom[067] = 8'h43; 
        rom[068] = 8'h44; 
        rom[069] = 8'h45; 
        rom[070] = 8'h46; 
        rom[071] = 8'h47; 
        rom[072] = 8'h48; 
        rom[073] = 8'h49; 
        rom[074] = 8'h4a; 
        rom[075] = 8'h4b; 
        rom[076] = 8'h4c; 
        rom[077] = 8'h4d; 
        rom[078] = 8'h4e; 
        rom[079] = 8'h4f; 
        rom[080] = 8'h50; 
        rom[081] = 8'h51; 
        rom[082] = 8'h52; 
        rom[083] = 8'h53; 
        rom[084] = 8'h54; 
        rom[085] = 8'h55; 
        rom[086] = 8'h56; 
        rom[087] = 8'h57; 
        rom[088] = 8'h58; 
        rom[089] = 8'h59; 
        rom[090] = 8'h5a; 
        rom[091] = 8'h5b; 
        rom[092] = 8'h5c; 
        rom[093] = 8'h5d; 
        rom[094] = 8'h5e; 
        rom[095] = 8'h5f; 
        rom[096] = 8'h60; 
        rom[097] = 8'h61; 
        rom[098] = 8'h62; 
        rom[099] = 8'h63; 
        rom[100] = 8'h64; 
        rom[101] = 8'h65; 
        rom[102] = 8'h66; 
        rom[103] = 8'h67; 
        rom[104] = 8'h68; 
        rom[105] = 8'h69; 
        rom[106] = 8'h6a; 
        rom[107] = 8'h6b; 
        rom[108] = 8'h6c; 
        rom[109] = 8'h6d; 
        rom[110] = 8'h6e; 
        rom[111] = 8'h6f; 
        rom[112] = 8'h70; 
        rom[113] = 8'h71; 
        rom[114] = 8'h72; 
        rom[115] = 8'h73; 
        rom[116] = 8'h74; 
        rom[117] = 8'h75; 
        rom[118] = 8'h76; 
        rom[119] = 8'h77; 
        rom[120] = 8'h78; 
        rom[121] = 8'h79; 
        rom[122] = 8'h7a; 
        rom[123] = 8'h7b; 
        rom[124] = 8'h7c; 
        rom[125] = 8'h7d; 
        rom[126] = 8'h7e; 
        rom[127] = 8'h7f; 
        rom[128] = 8'h80; 
        rom[129] = 8'h81; 
        rom[130] = 8'h82; 
        rom[131] = 8'h83; 
        rom[132] = 8'h84; 
        rom[133] = 8'h85; 
        rom[134] = 8'h86; 
        rom[135] = 8'h87; 
        rom[136] = 8'h88; 
        rom[137] = 8'h89; 
        rom[138] = 8'h8a; 
        rom[139] = 8'h8b; 
        rom[140] = 8'h8c; 
        rom[141] = 8'h8d; 
        rom[142] = 8'h8e; 
        rom[143] = 8'h8f; 
        rom[144] = 8'h90; 
        rom[145] = 8'h91; 
        rom[146] = 8'h92; 
        rom[147] = 8'h93; 
        rom[148] = 8'h94; 
        rom[149] = 8'h95; 
        rom[150] = 8'h96; 
        rom[151] = 8'h97; 
        rom[152] = 8'h98; 
        rom[153] = 8'h99; 
        rom[154] = 8'h9a; 
        rom[155] = 8'h9b; 
        rom[156] = 8'h9c; 
        rom[157] = 8'h9d; 
        rom[158] = 8'h9e; 
        rom[159] = 8'h9f; 
        rom[160] = 8'ha0; 
        rom[161] = 8'ha1; 
        rom[162] = 8'ha2; 
        rom[163] = 8'ha3; 
        rom[164] = 8'ha4; 
        rom[165] = 8'ha5; 
        rom[166] = 8'ha6; 
        rom[167] = 8'ha7; 
        rom[168] = 8'ha8; 
        rom[169] = 8'ha9; 
        rom[170] = 8'haa; 
        rom[171] = 8'hab; 
        rom[172] = 8'hac; 
        rom[173] = 8'had; 
        rom[174] = 8'hae; 
        rom[175] = 8'haf; 
        rom[176] = 8'hb0; 
        rom[177] = 8'hb1; 
        rom[178] = 8'hb2; 
        rom[179] = 8'hb3; 
        rom[180] = 8'hb4; 
        rom[181] = 8'hb5; 
        rom[182] = 8'hb6; 
        rom[183] = 8'hb7; 
        rom[184] = 8'hb8; 
        rom[185] = 8'hb9; 
        rom[186] = 8'hba; 
        rom[187] = 8'hbb; 
        rom[188] = 8'hbc; 
        rom[189] = 8'hbd; 
        rom[190] = 8'hbe; 
        rom[191] = 8'hbf; 
        rom[192] = 8'hc0; 
        rom[193] = 8'hc1; 
        rom[194] = 8'hc2; 
        rom[195] = 8'hc3; 
        rom[196] = 8'hc4; 
        rom[197] = 8'hc5; 
        rom[198] = 8'hc6; 
        rom[199] = 8'hc7; 
        rom[200] = 8'hc8; 
        rom[201] = 8'hc9; 
        rom[202] = 8'hca; 
        rom[203] = 8'hcb; 
        rom[204] = 8'hcc; 
        rom[205] = 8'hcd; 
        rom[206] = 8'hce; 
        rom[207] = 8'hcf; 
        rom[208] = 8'hd0; 
        rom[209] = 8'hd1; 
        rom[210] = 8'hd2; 
        rom[211] = 8'hd3; 
        rom[212] = 8'hd4; 
        rom[213] = 8'hd5; 
        rom[214] = 8'hd6; 
        rom[215] = 8'hd7; 
        rom[216] = 8'hd8; 
        rom[217] = 8'hd9; 
        rom[218] = 8'hda; 
        rom[219] = 8'hdb; 
        rom[220] = 8'hdc; 
        rom[221] = 8'hdd; 
        rom[222] = 8'hde; 
        rom[223] = 8'hdf; 
        rom[224] = 8'he0; 
        rom[225] = 8'he1; 
        rom[226] = 8'he2; 
        rom[227] = 8'he3; 
        rom[228] = 8'he4; 
        rom[229] = 8'he5; 
        rom[230] = 8'he6; 
        rom[231] = 8'he7; 
        rom[232] = 8'he8; 
        rom[233] = 8'he9; 
        rom[234] = 8'hea; 
        rom[235] = 8'heb; 
        rom[236] = 8'hec; 
        rom[237] = 8'hed; 
        rom[238] = 8'hee; 
        rom[239] = 8'hef; 
        rom[240] = 8'hf0; 
        rom[241] = 8'hf1; 
        rom[242] = 8'hf2; 
        rom[243] = 8'hf3; 
        rom[244] = 8'hf4; 
        rom[245] = 8'hf5; 
        rom[246] = 8'hf6; 
        rom[247] = 8'hf7; 
        rom[248] = 8'hf8; 
        rom[249] = 8'hf9; 
        rom[250] = 8'hfa; 
        rom[251] = 8'hfb; 
        rom[252] = 8'hfc; 
        rom[253] = 8'hfd; 
        rom[254] = 8'hfe; 
        rom[255] = 8'hff;
    end

    always @ (posedge clk)
    begin
        q <= rom[addr];
    end

endmodule
